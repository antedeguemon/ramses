library verilog;
use verilog.vl_types.all;
entity Ramses_vlg_vec_tst is
end Ramses_vlg_vec_tst;
